library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;



package project_pkg is




end package;
	
package body project_pkg is
	
end package body project_pkg;