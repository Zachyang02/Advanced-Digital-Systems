library ads;
use ads.ads_fixed.all;
use ads.ads_complex_pkg.all;

package seed_table is 
	type seed_rom_type is array (natural range<>) of ads_complex;
	constant seed_rom:	seed_rom_type := (
		( re => to_ads_sfixed(-1.50000), im => to_ads_sfixed( 0.00000) ),
			( re => to_ads_sfixed(-1.49849), im => to_ads_sfixed( 0.04487) ),
			( re => to_ads_sfixed(-1.49396), im => to_ads_sfixed( 0.08971) ),
			( re => to_ads_sfixed(-1.48642), im => to_ads_sfixed( 0.13446) ),
			( re => to_ads_sfixed(-1.47589), im => to_ads_sfixed( 0.17909) ),
			( re => to_ads_sfixed(-1.46239), im => to_ads_sfixed( 0.22356) ),
			( re => to_ads_sfixed(-1.44594), im => to_ads_sfixed( 0.26784) ),
			( re => to_ads_sfixed(-1.42658), im => to_ads_sfixed( 0.31187) ),
			( re => to_ads_sfixed(-1.40435), im => to_ads_sfixed( 0.35562) ),
			( re => to_ads_sfixed(-1.37929), im => to_ads_sfixed( 0.39906) ),
			( re => to_ads_sfixed(-1.35145), im => to_ads_sfixed( 0.44213) ),
			( re => to_ads_sfixed(-1.32089), im => to_ads_sfixed( 0.48481) ),
			( re => to_ads_sfixed(-1.28767), im => to_ads_sfixed( 0.52706) ),
			( re => to_ads_sfixed(-1.25186), im => to_ads_sfixed( 0.56884) ),
			( re => to_ads_sfixed(-1.21353), im => to_ads_sfixed( 0.61010) ),
			( re => to_ads_sfixed(-1.17275), im => to_ads_sfixed( 0.65083) ),
			( re => to_ads_sfixed(-1.12961), im => to_ads_sfixed( 0.69096) ),
			( re => to_ads_sfixed(-1.08419), im => to_ads_sfixed( 0.73048) ),
			( re => to_ads_sfixed(-1.03659), im => to_ads_sfixed( 0.76935) ),
			( re => to_ads_sfixed(-0.98691), im => to_ads_sfixed( 0.80753) ),
			( re => to_ads_sfixed(-0.93523), im => to_ads_sfixed( 0.84498) ),
			( re => to_ads_sfixed(-0.88168), im => to_ads_sfixed( 0.88168) ),
			( re => to_ads_sfixed(-0.82635), im => to_ads_sfixed( 0.91759) ),
			( re => to_ads_sfixed(-0.76935), im => to_ads_sfixed( 0.95267) ),
			( re => to_ads_sfixed(-0.71080), im => to_ads_sfixed( 0.98691) ),
			( re => to_ads_sfixed(-0.65083), im => to_ads_sfixed( 1.02026) ),
			( re => to_ads_sfixed(-0.58954), im => to_ads_sfixed( 1.05270) ),
			( re => to_ads_sfixed(-0.52706), im => to_ads_sfixed( 1.08419) ),
			( re => to_ads_sfixed(-0.46353), im => to_ads_sfixed( 1.11472) ),
			( re => to_ads_sfixed(-0.39906), im => to_ads_sfixed( 1.14424) ),
			( re => to_ads_sfixed(-0.33378), im => to_ads_sfixed( 1.17275) ),
			( re => to_ads_sfixed(-0.26784), im => to_ads_sfixed( 1.20020) ),
			( re => to_ads_sfixed(-0.20135), im => to_ads_sfixed( 1.22658) ),
			( re => to_ads_sfixed(-0.13446), im => to_ads_sfixed( 1.25186) ),
			( re => to_ads_sfixed(-0.06730), im => to_ads_sfixed( 1.27602) ),
			( re => to_ads_sfixed( 0.00000), im => to_ads_sfixed( 1.29904) ),
			( re => to_ads_sfixed( 0.06730), im => to_ads_sfixed( 1.32089) ),
			( re => to_ads_sfixed( 0.13446), im => to_ads_sfixed( 1.34157) ),
			( re => to_ads_sfixed( 0.20135), im => to_ads_sfixed( 1.36104) ),
			( re => to_ads_sfixed( 0.26784), im => to_ads_sfixed( 1.37929) ),
			( re => to_ads_sfixed( 0.33378), im => to_ads_sfixed( 1.39631) ),
			( re => to_ads_sfixed( 0.39906), im => to_ads_sfixed( 1.41208) ),
			( re => to_ads_sfixed( 0.46353), im => to_ads_sfixed( 1.42658) ),
			( re => to_ads_sfixed( 0.52706), im => to_ads_sfixed( 1.43981) ),
			( re => to_ads_sfixed( 0.58954), im => to_ads_sfixed( 1.45175) ),
			( re => to_ads_sfixed( 0.65083), im => to_ads_sfixed( 1.46239) ),
			( re => to_ads_sfixed( 0.71080), im => to_ads_sfixed( 1.47172) ),
			( re => to_ads_sfixed( 0.76935), im => to_ads_sfixed( 1.47974) ),
			( re => to_ads_sfixed( 0.82635), im => to_ads_sfixed( 1.48642) ),
			( re => to_ads_sfixed( 0.88168), im => to_ads_sfixed( 1.49178) ),
			( re => to_ads_sfixed( 0.93523), im => to_ads_sfixed( 1.49581) ),
			( re => to_ads_sfixed( 0.98691), im => to_ads_sfixed( 1.49849) ),
			( re => to_ads_sfixed( 1.03659), im => to_ads_sfixed( 1.49983) ),
			( re => to_ads_sfixed( 1.08419), im => to_ads_sfixed( 1.49983) ),
			( re => to_ads_sfixed( 1.12961), im => to_ads_sfixed( 1.49849) ),
			( re => to_ads_sfixed( 1.17275), im => to_ads_sfixed( 1.49581) ),
			( re => to_ads_sfixed( 1.21353), im => to_ads_sfixed( 1.49178) ),
			( re => to_ads_sfixed( 1.25186), im => to_ads_sfixed( 1.48642) ),
			( re => to_ads_sfixed( 1.28767), im => to_ads_sfixed( 1.47974) ),
			( re => to_ads_sfixed( 1.32089), im => to_ads_sfixed( 1.47172) ),
			( re => to_ads_sfixed( 1.35145), im => to_ads_sfixed( 1.46239) ),
			( re => to_ads_sfixed( 1.37929), im => to_ads_sfixed( 1.45175) ),
			( re => to_ads_sfixed( 1.40435), im => to_ads_sfixed( 1.43981) ),
			( re => to_ads_sfixed( 1.42658), im => to_ads_sfixed( 1.42658) ),
			( re => to_ads_sfixed( 1.44594), im => to_ads_sfixed( 1.41208) ),
			( re => to_ads_sfixed( 1.46239), im => to_ads_sfixed( 1.39631) ),
			( re => to_ads_sfixed( 1.47589), im => to_ads_sfixed( 1.37929) ),
			( re => to_ads_sfixed( 1.48642), im => to_ads_sfixed( 1.36104) ),
			( re => to_ads_sfixed( 1.49396), im => to_ads_sfixed( 1.34157) ),
			( re => to_ads_sfixed( 1.49849), im => to_ads_sfixed( 1.32089) ),
			( re => to_ads_sfixed( 1.50000), im => to_ads_sfixed( 1.29904) ),
			( re => to_ads_sfixed( 1.49849), im => to_ads_sfixed( 1.27602) ),
			( re => to_ads_sfixed( 1.49396), im => to_ads_sfixed( 1.25186) ),
			( re => to_ads_sfixed( 1.48642), im => to_ads_sfixed( 1.22658) ),
			( re => to_ads_sfixed( 1.47589), im => to_ads_sfixed( 1.20020) ),
			( re => to_ads_sfixed( 1.46239), im => to_ads_sfixed( 1.17275) ),
			( re => to_ads_sfixed( 1.44594), im => to_ads_sfixed( 1.14424) ),
			( re => to_ads_sfixed( 1.42658), im => to_ads_sfixed( 1.11472) ),
			( re => to_ads_sfixed( 1.40435), im => to_ads_sfixed( 1.08419) ),
			( re => to_ads_sfixed( 1.37929), im => to_ads_sfixed( 1.05270) ),
			( re => to_ads_sfixed( 1.35145), im => to_ads_sfixed( 1.02026) ),
			( re => to_ads_sfixed( 1.32089), im => to_ads_sfixed( 0.98691) ),
			( re => to_ads_sfixed( 1.28767), im => to_ads_sfixed( 0.95267) ),
			( re => to_ads_sfixed( 1.25186), im => to_ads_sfixed( 0.91759) ),
			( re => to_ads_sfixed( 1.21353), im => to_ads_sfixed( 0.88168) ),
			( re => to_ads_sfixed( 1.17275), im => to_ads_sfixed( 0.84498) ),
			( re => to_ads_sfixed( 1.12961), im => to_ads_sfixed( 0.80753) ),
			( re => to_ads_sfixed( 1.08419), im => to_ads_sfixed( 0.76935) ),
			( re => to_ads_sfixed( 1.03659), im => to_ads_sfixed( 0.73048) ),
			( re => to_ads_sfixed( 0.98691), im => to_ads_sfixed( 0.69096) ),
			( re => to_ads_sfixed( 0.93523), im => to_ads_sfixed( 0.65083) ),
			( re => to_ads_sfixed( 0.88168), im => to_ads_sfixed( 0.61010) ),
			( re => to_ads_sfixed( 0.82635), im => to_ads_sfixed( 0.56884) ),
			( re => to_ads_sfixed( 0.76935), im => to_ads_sfixed( 0.52706) ),
			( re => to_ads_sfixed( 0.71080), im => to_ads_sfixed( 0.48481) ),
			( re => to_ads_sfixed( 0.65083), im => to_ads_sfixed( 0.44213) ),
			( re => to_ads_sfixed( 0.58954), im => to_ads_sfixed( 0.39906) ),
			( re => to_ads_sfixed( 0.52706), im => to_ads_sfixed( 0.35562) ),
			( re => to_ads_sfixed( 0.46353), im => to_ads_sfixed( 0.31187) ),
			( re => to_ads_sfixed( 0.39906), im => to_ads_sfixed( 0.26784) ),
			( re => to_ads_sfixed( 0.33378), im => to_ads_sfixed( 0.22356) ),
			( re => to_ads_sfixed( 0.26784), im => to_ads_sfixed( 0.17909) ),
			( re => to_ads_sfixed( 0.20135), im => to_ads_sfixed( 0.13446) ),
			( re => to_ads_sfixed( 0.13446), im => to_ads_sfixed( 0.08971) ),
			( re => to_ads_sfixed( 0.06730), im => to_ads_sfixed( 0.04487) ),
			( re => to_ads_sfixed(-0.00000), im => to_ads_sfixed(-0.00000) ),
			( re => to_ads_sfixed(-0.06730), im => to_ads_sfixed(-0.04487) ),
			( re => to_ads_sfixed(-0.13446), im => to_ads_sfixed(-0.08971) ),
			( re => to_ads_sfixed(-0.20135), im => to_ads_sfixed(-0.13446) ),
			( re => to_ads_sfixed(-0.26784), im => to_ads_sfixed(-0.17909) ),
			( re => to_ads_sfixed(-0.33378), im => to_ads_sfixed(-0.22356) ),
			( re => to_ads_sfixed(-0.39906), im => to_ads_sfixed(-0.26784) ),
			( re => to_ads_sfixed(-0.46353), im => to_ads_sfixed(-0.31187) ),
			( re => to_ads_sfixed(-0.52706), im => to_ads_sfixed(-0.35562) ),
			( re => to_ads_sfixed(-0.58954), im => to_ads_sfixed(-0.39906) ),
			( re => to_ads_sfixed(-0.65083), im => to_ads_sfixed(-0.44213) ),
			( re => to_ads_sfixed(-0.71080), im => to_ads_sfixed(-0.48481) ),
			( re => to_ads_sfixed(-0.76935), im => to_ads_sfixed(-0.52706) ),
			( re => to_ads_sfixed(-0.82635), im => to_ads_sfixed(-0.56884) ),
			( re => to_ads_sfixed(-0.88168), im => to_ads_sfixed(-0.61010) ),
			( re => to_ads_sfixed(-0.93523), im => to_ads_sfixed(-0.65083) ),
			( re => to_ads_sfixed(-0.98691), im => to_ads_sfixed(-0.69096) ),
			( re => to_ads_sfixed(-1.03659), im => to_ads_sfixed(-0.73048) ),
			( re => to_ads_sfixed(-1.08419), im => to_ads_sfixed(-0.76935) ),
			( re => to_ads_sfixed(-1.12961), im => to_ads_sfixed(-0.80753) ),
			( re => to_ads_sfixed(-1.17275), im => to_ads_sfixed(-0.84498) ),
			( re => to_ads_sfixed(-1.21353), im => to_ads_sfixed(-0.88168) ),
			( re => to_ads_sfixed(-1.25186), im => to_ads_sfixed(-0.91759) ),
			( re => to_ads_sfixed(-1.28767), im => to_ads_sfixed(-0.95267) ),
			( re => to_ads_sfixed(-1.32089), im => to_ads_sfixed(-0.98691) ),
			( re => to_ads_sfixed(-1.35145), im => to_ads_sfixed(-1.02026) ),
			( re => to_ads_sfixed(-1.37929), im => to_ads_sfixed(-1.05270) ),
			( re => to_ads_sfixed(-1.40435), im => to_ads_sfixed(-1.08419) ),
			( re => to_ads_sfixed(-1.42658), im => to_ads_sfixed(-1.11472) ),
			( re => to_ads_sfixed(-1.44594), im => to_ads_sfixed(-1.14424) ),
			( re => to_ads_sfixed(-1.46239), im => to_ads_sfixed(-1.17275) ),
			( re => to_ads_sfixed(-1.47589), im => to_ads_sfixed(-1.20020) ),
			( re => to_ads_sfixed(-1.48642), im => to_ads_sfixed(-1.22658) ),
			( re => to_ads_sfixed(-1.49396), im => to_ads_sfixed(-1.25186) ),
			( re => to_ads_sfixed(-1.49849), im => to_ads_sfixed(-1.27602) ),
			( re => to_ads_sfixed(-1.50000), im => to_ads_sfixed(-1.29904) ),
			( re => to_ads_sfixed(-1.49849), im => to_ads_sfixed(-1.32089) ),
			( re => to_ads_sfixed(-1.49396), im => to_ads_sfixed(-1.34157) ),
			( re => to_ads_sfixed(-1.48642), im => to_ads_sfixed(-1.36104) ),
			( re => to_ads_sfixed(-1.47589), im => to_ads_sfixed(-1.37929) ),
			( re => to_ads_sfixed(-1.46239), im => to_ads_sfixed(-1.39631) ),
			( re => to_ads_sfixed(-1.44594), im => to_ads_sfixed(-1.41208) ),
			( re => to_ads_sfixed(-1.42658), im => to_ads_sfixed(-1.42658) ),
			( re => to_ads_sfixed(-1.40435), im => to_ads_sfixed(-1.43981) ),
			( re => to_ads_sfixed(-1.37929), im => to_ads_sfixed(-1.45175) ),
			( re => to_ads_sfixed(-1.35145), im => to_ads_sfixed(-1.46239) ),
			( re => to_ads_sfixed(-1.32089), im => to_ads_sfixed(-1.47172) ),
			( re => to_ads_sfixed(-1.28767), im => to_ads_sfixed(-1.47974) ),
			( re => to_ads_sfixed(-1.25186), im => to_ads_sfixed(-1.48642) ),
			( re => to_ads_sfixed(-1.21353), im => to_ads_sfixed(-1.49178) ),
			( re => to_ads_sfixed(-1.17275), im => to_ads_sfixed(-1.49581) ),
			( re => to_ads_sfixed(-1.12961), im => to_ads_sfixed(-1.49849) ),
			( re => to_ads_sfixed(-1.08419), im => to_ads_sfixed(-1.49983) ),
			( re => to_ads_sfixed(-1.03659), im => to_ads_sfixed(-1.49983) ),
			( re => to_ads_sfixed(-0.98691), im => to_ads_sfixed(-1.49849) ),
			( re => to_ads_sfixed(-0.93523), im => to_ads_sfixed(-1.49581) ),
			( re => to_ads_sfixed(-0.88168), im => to_ads_sfixed(-1.49178) ),
			( re => to_ads_sfixed(-0.82635), im => to_ads_sfixed(-1.48642) ),
			( re => to_ads_sfixed(-0.76935), im => to_ads_sfixed(-1.47974) ),
			( re => to_ads_sfixed(-0.71080), im => to_ads_sfixed(-1.47172) ),
			( re => to_ads_sfixed(-0.65083), im => to_ads_sfixed(-1.46239) ),
			( re => to_ads_sfixed(-0.58954), im => to_ads_sfixed(-1.45175) ),
			( re => to_ads_sfixed(-0.52706), im => to_ads_sfixed(-1.43981) ),
			( re => to_ads_sfixed(-0.46353), im => to_ads_sfixed(-1.42658) ),
			( re => to_ads_sfixed(-0.39906), im => to_ads_sfixed(-1.41208) ),
			( re => to_ads_sfixed(-0.33378), im => to_ads_sfixed(-1.39631) ),
			( re => to_ads_sfixed(-0.26784), im => to_ads_sfixed(-1.37929) ),
			( re => to_ads_sfixed(-0.20135), im => to_ads_sfixed(-1.36104) ),
			( re => to_ads_sfixed(-0.13446), im => to_ads_sfixed(-1.34157) ),
			( re => to_ads_sfixed(-0.06730), im => to_ads_sfixed(-1.32089) ),
			( re => to_ads_sfixed( 0.00000), im => to_ads_sfixed(-1.29904) ),
			( re => to_ads_sfixed( 0.06730), im => to_ads_sfixed(-1.27602) ),
			( re => to_ads_sfixed( 0.13446), im => to_ads_sfixed(-1.25186) ),
			( re => to_ads_sfixed( 0.20135), im => to_ads_sfixed(-1.22658) ),
			( re => to_ads_sfixed( 0.26784), im => to_ads_sfixed(-1.20020) ),
			( re => to_ads_sfixed( 0.33378), im => to_ads_sfixed(-1.17275) ),
			( re => to_ads_sfixed( 0.39906), im => to_ads_sfixed(-1.14424) ),
			( re => to_ads_sfixed( 0.46353), im => to_ads_sfixed(-1.11472) ),
			( re => to_ads_sfixed( 0.52706), im => to_ads_sfixed(-1.08419) ),
			( re => to_ads_sfixed( 0.58954), im => to_ads_sfixed(-1.05270) ),
			( re => to_ads_sfixed( 0.65083), im => to_ads_sfixed(-1.02026) ),
			( re => to_ads_sfixed( 0.71080), im => to_ads_sfixed(-0.98691) ),
			( re => to_ads_sfixed( 0.76935), im => to_ads_sfixed(-0.95267) ),
			( re => to_ads_sfixed( 0.82635), im => to_ads_sfixed(-0.91759) ),
			( re => to_ads_sfixed( 0.88168), im => to_ads_sfixed(-0.88168) ),
			( re => to_ads_sfixed( 0.93523), im => to_ads_sfixed(-0.84498) ),
			( re => to_ads_sfixed( 0.98691), im => to_ads_sfixed(-0.80753) ),
			( re => to_ads_sfixed( 1.03659), im => to_ads_sfixed(-0.76935) ),
			( re => to_ads_sfixed( 1.08419), im => to_ads_sfixed(-0.73048) ),
			( re => to_ads_sfixed( 1.12961), im => to_ads_sfixed(-0.69096) ),
			( re => to_ads_sfixed( 1.17275), im => to_ads_sfixed(-0.65083) ),
			( re => to_ads_sfixed( 1.21353), im => to_ads_sfixed(-0.61010) ),
			( re => to_ads_sfixed( 1.25186), im => to_ads_sfixed(-0.56884) ),
			( re => to_ads_sfixed( 1.28767), im => to_ads_sfixed(-0.52706) ),
			( re => to_ads_sfixed( 1.32089), im => to_ads_sfixed(-0.48481) ),
			( re => to_ads_sfixed( 1.35145), im => to_ads_sfixed(-0.44213) ),
			( re => to_ads_sfixed( 1.37929), im => to_ads_sfixed(-0.39906) ),
			( re => to_ads_sfixed( 1.40435), im => to_ads_sfixed(-0.35562) ),
			( re => to_ads_sfixed( 1.42658), im => to_ads_sfixed(-0.31187) ),
			( re => to_ads_sfixed( 1.44594), im => to_ads_sfixed(-0.26784) ),
			( re => to_ads_sfixed( 1.46239), im => to_ads_sfixed(-0.22356) ),
			( re => to_ads_sfixed( 1.47589), im => to_ads_sfixed(-0.17909) ),
			( re => to_ads_sfixed( 1.48642), im => to_ads_sfixed(-0.13446) ),
			( re => to_ads_sfixed( 1.49396), im => to_ads_sfixed(-0.08971) ),
			( re => to_ads_sfixed( 1.49849), im => to_ads_sfixed(-0.04487) ),
			( re => to_ads_sfixed( 1.50000), im => to_ads_sfixed( 0.00000) ),
			( re => to_ads_sfixed( 1.49849), im => to_ads_sfixed( 0.04487) ),
			( re => to_ads_sfixed( 1.49396), im => to_ads_sfixed( 0.08971) ),
			( re => to_ads_sfixed( 1.48642), im => to_ads_sfixed( 0.13446) ),
			( re => to_ads_sfixed( 1.47589), im => to_ads_sfixed( 0.17909) ),
			( re => to_ads_sfixed( 1.46239), im => to_ads_sfixed( 0.22356) ),
			( re => to_ads_sfixed( 1.44594), im => to_ads_sfixed( 0.26784) ),
			( re => to_ads_sfixed( 1.42658), im => to_ads_sfixed( 0.31187) ),
			( re => to_ads_sfixed( 1.40435), im => to_ads_sfixed( 0.35562) ),
			( re => to_ads_sfixed( 1.37929), im => to_ads_sfixed( 0.39906) ),
			( re => to_ads_sfixed( 1.35145), im => to_ads_sfixed( 0.44213) ),
			( re => to_ads_sfixed( 1.32089), im => to_ads_sfixed( 0.48481) ),
			( re => to_ads_sfixed( 1.28767), im => to_ads_sfixed( 0.52706) ),
			( re => to_ads_sfixed( 1.25186), im => to_ads_sfixed( 0.56884) ),
			( re => to_ads_sfixed( 1.21353), im => to_ads_sfixed( 0.61010) ),
			( re => to_ads_sfixed( 1.17275), im => to_ads_sfixed( 0.65083) ),
			( re => to_ads_sfixed( 1.12961), im => to_ads_sfixed( 0.69096) ),
			( re => to_ads_sfixed( 1.08419), im => to_ads_sfixed( 0.73048) ),
			( re => to_ads_sfixed( 1.03659), im => to_ads_sfixed( 0.76935) ),
			( re => to_ads_sfixed( 0.98691), im => to_ads_sfixed( 0.80753) ),
			( re => to_ads_sfixed( 0.93523), im => to_ads_sfixed( 0.84498) ),
			( re => to_ads_sfixed( 0.88168), im => to_ads_sfixed( 0.88168) ),
			( re => to_ads_sfixed( 0.82635), im => to_ads_sfixed( 0.91759) ),
			( re => to_ads_sfixed( 0.76935), im => to_ads_sfixed( 0.95267) ),
			( re => to_ads_sfixed( 0.71080), im => to_ads_sfixed( 0.98691) ),
			( re => to_ads_sfixed( 0.65083), im => to_ads_sfixed( 1.02026) ),
			( re => to_ads_sfixed( 0.58954), im => to_ads_sfixed( 1.05270) ),
			( re => to_ads_sfixed( 0.52706), im => to_ads_sfixed( 1.08419) ),
			( re => to_ads_sfixed( 0.46353), im => to_ads_sfixed( 1.11472) ),
			( re => to_ads_sfixed( 0.39906), im => to_ads_sfixed( 1.14424) ),
			( re => to_ads_sfixed( 0.33378), im => to_ads_sfixed( 1.17275) ),
			( re => to_ads_sfixed( 0.26784), im => to_ads_sfixed( 1.20020) ),
			( re => to_ads_sfixed( 0.20135), im => to_ads_sfixed( 1.22658) ),
			( re => to_ads_sfixed( 0.13446), im => to_ads_sfixed( 1.25186) ),
			( re => to_ads_sfixed( 0.06730), im => to_ads_sfixed( 1.27602) ),
			( re => to_ads_sfixed(-0.00000), im => to_ads_sfixed( 1.29904) ),
			( re => to_ads_sfixed(-0.06730), im => to_ads_sfixed( 1.32089) ),
			( re => to_ads_sfixed(-0.13446), im => to_ads_sfixed( 1.34157) ),
			( re => to_ads_sfixed(-0.20135), im => to_ads_sfixed( 1.36104) ),
			( re => to_ads_sfixed(-0.26784), im => to_ads_sfixed( 1.37929) ),
			( re => to_ads_sfixed(-0.33378), im => to_ads_sfixed( 1.39631) ),
			( re => to_ads_sfixed(-0.39906), im => to_ads_sfixed( 1.41208) ),
			( re => to_ads_sfixed(-0.46353), im => to_ads_sfixed( 1.42658) ),
			( re => to_ads_sfixed(-0.52706), im => to_ads_sfixed( 1.43981) ),
			( re => to_ads_sfixed(-0.58954), im => to_ads_sfixed( 1.45175) ),
			( re => to_ads_sfixed(-0.65083), im => to_ads_sfixed( 1.46239) ),
			( re => to_ads_sfixed(-0.71080), im => to_ads_sfixed( 1.47172) ),
			( re => to_ads_sfixed(-0.76935), im => to_ads_sfixed( 1.47974) ),
			( re => to_ads_sfixed(-0.82635), im => to_ads_sfixed( 1.48642) ),
			( re => to_ads_sfixed(-0.88168), im => to_ads_sfixed( 1.49178) ),
			( re => to_ads_sfixed(-0.93523), im => to_ads_sfixed( 1.49581) ),
			( re => to_ads_sfixed(-0.98691), im => to_ads_sfixed( 1.49849) ),
			( re => to_ads_sfixed(-1.03659), im => to_ads_sfixed( 1.49983) ),
			( re => to_ads_sfixed(-1.08419), im => to_ads_sfixed( 1.49983) ),
			( re => to_ads_sfixed(-1.12961), im => to_ads_sfixed( 1.49849) ),
			( re => to_ads_sfixed(-1.17275), im => to_ads_sfixed( 1.49581) ),
			( re => to_ads_sfixed(-1.21353), im => to_ads_sfixed( 1.49178) ),
			( re => to_ads_sfixed(-1.25186), im => to_ads_sfixed( 1.48642) ),
			( re => to_ads_sfixed(-1.28767), im => to_ads_sfixed( 1.47974) ),
			( re => to_ads_sfixed(-1.32089), im => to_ads_sfixed( 1.47172) ),
			( re => to_ads_sfixed(-1.35145), im => to_ads_sfixed( 1.46239) ),
			( re => to_ads_sfixed(-1.37929), im => to_ads_sfixed( 1.45175) ),
			( re => to_ads_sfixed(-1.40435), im => to_ads_sfixed( 1.43981) ),
			( re => to_ads_sfixed(-1.42658), im => to_ads_sfixed( 1.42658) ),
			( re => to_ads_sfixed(-1.44594), im => to_ads_sfixed( 1.41208) ),
			( re => to_ads_sfixed(-1.46239), im => to_ads_sfixed( 1.39631) ),
			( re => to_ads_sfixed(-1.47589), im => to_ads_sfixed( 1.37929) ),
			( re => to_ads_sfixed(-1.48642), im => to_ads_sfixed( 1.36104) ),
			( re => to_ads_sfixed(-1.49396), im => to_ads_sfixed( 1.34157) ),
			( re => to_ads_sfixed(-1.49849), im => to_ads_sfixed( 1.32089) ),
			( re => to_ads_sfixed(-1.50000), im => to_ads_sfixed( 1.29904) ),
			( re => to_ads_sfixed(-1.49849), im => to_ads_sfixed( 1.27602) ),
			( re => to_ads_sfixed(-1.49396), im => to_ads_sfixed( 1.25186) ),
			( re => to_ads_sfixed(-1.48642), im => to_ads_sfixed( 1.22658) ),
			( re => to_ads_sfixed(-1.47589), im => to_ads_sfixed( 1.20020) ),
			( re => to_ads_sfixed(-1.46239), im => to_ads_sfixed( 1.17275) ),
			( re => to_ads_sfixed(-1.44594), im => to_ads_sfixed( 1.14424) ),
			( re => to_ads_sfixed(-1.42658), im => to_ads_sfixed( 1.11472) ),
			( re => to_ads_sfixed(-1.40435), im => to_ads_sfixed( 1.08419) ),
			( re => to_ads_sfixed(-1.37929), im => to_ads_sfixed( 1.05270) ),
			( re => to_ads_sfixed(-1.35145), im => to_ads_sfixed( 1.02026) ),
			( re => to_ads_sfixed(-1.32089), im => to_ads_sfixed( 0.98691) ),
			( re => to_ads_sfixed(-1.28767), im => to_ads_sfixed( 0.95267) ),
			( re => to_ads_sfixed(-1.25186), im => to_ads_sfixed( 0.91759) ),
			( re => to_ads_sfixed(-1.21353), im => to_ads_sfixed( 0.88168) ),
			( re => to_ads_sfixed(-1.17275), im => to_ads_sfixed( 0.84498) ),
			( re => to_ads_sfixed(-1.12961), im => to_ads_sfixed( 0.80753) ),
			( re => to_ads_sfixed(-1.08419), im => to_ads_sfixed( 0.76935) ),
			( re => to_ads_sfixed(-1.03659), im => to_ads_sfixed( 0.73048) ),
			( re => to_ads_sfixed(-0.98691), im => to_ads_sfixed( 0.69096) ),
			( re => to_ads_sfixed(-0.93523), im => to_ads_sfixed( 0.65083) ),
			( re => to_ads_sfixed(-0.88168), im => to_ads_sfixed( 0.61010) ),
			( re => to_ads_sfixed(-0.82635), im => to_ads_sfixed( 0.56884) ),
			( re => to_ads_sfixed(-0.76935), im => to_ads_sfixed( 0.52706) ),
			( re => to_ads_sfixed(-0.71080), im => to_ads_sfixed( 0.48481) ),
			( re => to_ads_sfixed(-0.65083), im => to_ads_sfixed( 0.44213) ),
			( re => to_ads_sfixed(-0.58954), im => to_ads_sfixed( 0.39906) ),
			( re => to_ads_sfixed(-0.52706), im => to_ads_sfixed( 0.35562) ),
			( re => to_ads_sfixed(-0.46353), im => to_ads_sfixed( 0.31187) ),
			( re => to_ads_sfixed(-0.39906), im => to_ads_sfixed( 0.26784) ),
			( re => to_ads_sfixed(-0.33378), im => to_ads_sfixed( 0.22356) ),
			( re => to_ads_sfixed(-0.26784), im => to_ads_sfixed( 0.17909) ),
			( re => to_ads_sfixed(-0.20135), im => to_ads_sfixed( 0.13446) ),
			( re => to_ads_sfixed(-0.13446), im => to_ads_sfixed( 0.08971) ),
			( re => to_ads_sfixed(-0.06730), im => to_ads_sfixed( 0.04487) ),
			( re => to_ads_sfixed(-0.00000), im => to_ads_sfixed( 0.00000) ),
			( re => to_ads_sfixed( 0.06730), im => to_ads_sfixed(-0.04487) ),
			( re => to_ads_sfixed( 0.13446), im => to_ads_sfixed(-0.08971) ),
			( re => to_ads_sfixed( 0.20135), im => to_ads_sfixed(-0.13446) ),
			( re => to_ads_sfixed( 0.26784), im => to_ads_sfixed(-0.17909) ),
			( re => to_ads_sfixed( 0.33378), im => to_ads_sfixed(-0.22356) ),
			( re => to_ads_sfixed( 0.39906), im => to_ads_sfixed(-0.26784) ),
			( re => to_ads_sfixed( 0.46353), im => to_ads_sfixed(-0.31187) ),
			( re => to_ads_sfixed( 0.52706), im => to_ads_sfixed(-0.35562) ),
			( re => to_ads_sfixed( 0.58954), im => to_ads_sfixed(-0.39906) ),
			( re => to_ads_sfixed( 0.65083), im => to_ads_sfixed(-0.44213) ),
			( re => to_ads_sfixed( 0.71080), im => to_ads_sfixed(-0.48481) ),
			( re => to_ads_sfixed( 0.76935), im => to_ads_sfixed(-0.52706) ),
			( re => to_ads_sfixed( 0.82635), im => to_ads_sfixed(-0.56884) ),
			( re => to_ads_sfixed( 0.88168), im => to_ads_sfixed(-0.61010) ),
			( re => to_ads_sfixed( 0.93523), im => to_ads_sfixed(-0.65083) ),
			( re => to_ads_sfixed( 0.98691), im => to_ads_sfixed(-0.69096) ),
			( re => to_ads_sfixed( 1.03659), im => to_ads_sfixed(-0.73048) ),
			( re => to_ads_sfixed( 1.08419), im => to_ads_sfixed(-0.76935) ),
			( re => to_ads_sfixed( 1.12961), im => to_ads_sfixed(-0.80753) ),
			( re => to_ads_sfixed( 1.17275), im => to_ads_sfixed(-0.84498) ),
			( re => to_ads_sfixed( 1.21353), im => to_ads_sfixed(-0.88168) ),
			( re => to_ads_sfixed( 1.25186), im => to_ads_sfixed(-0.91759) ),
			( re => to_ads_sfixed( 1.28767), im => to_ads_sfixed(-0.95267) ),
			( re => to_ads_sfixed( 1.32089), im => to_ads_sfixed(-0.98691) ),
			( re => to_ads_sfixed( 1.35145), im => to_ads_sfixed(-1.02026) ),
			( re => to_ads_sfixed( 1.37929), im => to_ads_sfixed(-1.05270) ),
			( re => to_ads_sfixed( 1.40435), im => to_ads_sfixed(-1.08419) ),
			( re => to_ads_sfixed( 1.42658), im => to_ads_sfixed(-1.11472) ),
			( re => to_ads_sfixed( 1.44594), im => to_ads_sfixed(-1.14424) ),
			( re => to_ads_sfixed( 1.46239), im => to_ads_sfixed(-1.17275) ),
			( re => to_ads_sfixed( 1.47589), im => to_ads_sfixed(-1.20020) ),
			( re => to_ads_sfixed( 1.48642), im => to_ads_sfixed(-1.22658) ),
			( re => to_ads_sfixed( 1.49396), im => to_ads_sfixed(-1.25186) ),
			( re => to_ads_sfixed( 1.49849), im => to_ads_sfixed(-1.27602) ),
			( re => to_ads_sfixed( 1.50000), im => to_ads_sfixed(-1.29904) ),
			( re => to_ads_sfixed( 1.49849), im => to_ads_sfixed(-1.32089) ),
			( re => to_ads_sfixed( 1.49396), im => to_ads_sfixed(-1.34157) ),
			( re => to_ads_sfixed( 1.48642), im => to_ads_sfixed(-1.36104) ),
			( re => to_ads_sfixed( 1.47589), im => to_ads_sfixed(-1.37929) ),
			( re => to_ads_sfixed( 1.46239), im => to_ads_sfixed(-1.39631) ),
			( re => to_ads_sfixed( 1.44594), im => to_ads_sfixed(-1.41208) ),
			( re => to_ads_sfixed( 1.42658), im => to_ads_sfixed(-1.42658) ),
			( re => to_ads_sfixed( 1.40435), im => to_ads_sfixed(-1.43981) ),
			( re => to_ads_sfixed( 1.37929), im => to_ads_sfixed(-1.45175) ),
			( re => to_ads_sfixed( 1.35145), im => to_ads_sfixed(-1.46239) ),
			( re => to_ads_sfixed( 1.32089), im => to_ads_sfixed(-1.47172) ),
			( re => to_ads_sfixed( 1.28767), im => to_ads_sfixed(-1.47974) ),
			( re => to_ads_sfixed( 1.25186), im => to_ads_sfixed(-1.48642) ),
			( re => to_ads_sfixed( 1.21353), im => to_ads_sfixed(-1.49178) ),
			( re => to_ads_sfixed( 1.17275), im => to_ads_sfixed(-1.49581) ),
			( re => to_ads_sfixed( 1.12961), im => to_ads_sfixed(-1.49849) ),
			( re => to_ads_sfixed( 1.08419), im => to_ads_sfixed(-1.49983) ),
			( re => to_ads_sfixed( 1.03659), im => to_ads_sfixed(-1.49983) ),
			( re => to_ads_sfixed( 0.98691), im => to_ads_sfixed(-1.49849) ),
			( re => to_ads_sfixed( 0.93523), im => to_ads_sfixed(-1.49581) ),
			( re => to_ads_sfixed( 0.88168), im => to_ads_sfixed(-1.49178) ),
			( re => to_ads_sfixed( 0.82635), im => to_ads_sfixed(-1.48642) ),
			( re => to_ads_sfixed( 0.76935), im => to_ads_sfixed(-1.47974) ),
			( re => to_ads_sfixed( 0.71080), im => to_ads_sfixed(-1.47172) ),
			( re => to_ads_sfixed( 0.65083), im => to_ads_sfixed(-1.46239) ),
			( re => to_ads_sfixed( 0.58954), im => to_ads_sfixed(-1.45175) ),
			( re => to_ads_sfixed( 0.52706), im => to_ads_sfixed(-1.43981) ),
			( re => to_ads_sfixed( 0.46353), im => to_ads_sfixed(-1.42658) ),
			( re => to_ads_sfixed( 0.39906), im => to_ads_sfixed(-1.41208) ),
			( re => to_ads_sfixed( 0.33378), im => to_ads_sfixed(-1.39631) ),
			( re => to_ads_sfixed( 0.26784), im => to_ads_sfixed(-1.37929) ),
			( re => to_ads_sfixed( 0.20135), im => to_ads_sfixed(-1.36104) ),
			( re => to_ads_sfixed( 0.13446), im => to_ads_sfixed(-1.34157) ),
			( re => to_ads_sfixed( 0.06730), im => to_ads_sfixed(-1.32089) ),
			( re => to_ads_sfixed(-0.00000), im => to_ads_sfixed(-1.29904) ),
			( re => to_ads_sfixed(-0.06730), im => to_ads_sfixed(-1.27602) ),
			( re => to_ads_sfixed(-0.13446), im => to_ads_sfixed(-1.25186) ),
			( re => to_ads_sfixed(-0.20135), im => to_ads_sfixed(-1.22658) ),
			( re => to_ads_sfixed(-0.26784), im => to_ads_sfixed(-1.20020) ),
			( re => to_ads_sfixed(-0.33378), im => to_ads_sfixed(-1.17275) ),
			( re => to_ads_sfixed(-0.39906), im => to_ads_sfixed(-1.14424) ),
			( re => to_ads_sfixed(-0.46353), im => to_ads_sfixed(-1.11472) ),
			( re => to_ads_sfixed(-0.52706), im => to_ads_sfixed(-1.08419) ),
			( re => to_ads_sfixed(-0.58954), im => to_ads_sfixed(-1.05270) ),
			( re => to_ads_sfixed(-0.65083), im => to_ads_sfixed(-1.02026) ),
			( re => to_ads_sfixed(-0.71080), im => to_ads_sfixed(-0.98691) ),
			( re => to_ads_sfixed(-0.76935), im => to_ads_sfixed(-0.95267) ),
			( re => to_ads_sfixed(-0.82635), im => to_ads_sfixed(-0.91759) ),
			( re => to_ads_sfixed(-0.88168), im => to_ads_sfixed(-0.88168) ),
			( re => to_ads_sfixed(-0.93523), im => to_ads_sfixed(-0.84498) ),
			( re => to_ads_sfixed(-0.98691), im => to_ads_sfixed(-0.80753) ),
			( re => to_ads_sfixed(-1.03659), im => to_ads_sfixed(-0.76935) ),
			( re => to_ads_sfixed(-1.08419), im => to_ads_sfixed(-0.73048) ),
			( re => to_ads_sfixed(-1.12961), im => to_ads_sfixed(-0.69096) ),
			( re => to_ads_sfixed(-1.17275), im => to_ads_sfixed(-0.65083) ),
			( re => to_ads_sfixed(-1.21353), im => to_ads_sfixed(-0.61010) ),
			( re => to_ads_sfixed(-1.25186), im => to_ads_sfixed(-0.56884) ),
			( re => to_ads_sfixed(-1.28767), im => to_ads_sfixed(-0.52706) ),
			( re => to_ads_sfixed(-1.32089), im => to_ads_sfixed(-0.48481) ),
			( re => to_ads_sfixed(-1.35145), im => to_ads_sfixed(-0.44213) ),
			( re => to_ads_sfixed(-1.37929), im => to_ads_sfixed(-0.39906) ),
			( re => to_ads_sfixed(-1.40435), im => to_ads_sfixed(-0.35562) ),
			( re => to_ads_sfixed(-1.42658), im => to_ads_sfixed(-0.31187) ),
			( re => to_ads_sfixed(-1.44594), im => to_ads_sfixed(-0.26784) ),
			( re => to_ads_sfixed(-1.46239), im => to_ads_sfixed(-0.22356) ),
			( re => to_ads_sfixed(-1.47589), im => to_ads_sfixed(-0.17909) ),
			( re => to_ads_sfixed(-1.48642), im => to_ads_sfixed(-0.13446) ),
			( re => to_ads_sfixed(-1.49396), im => to_ads_sfixed(-0.08971) ),
			( re => to_ads_sfixed(-1.49849), im => to_ads_sfixed(-0.04487) )
	);
	
	
	constant seed_rom_total: natural := seed_rom'length;
	
	
	subtype seed_index_type is natural range 0 to seed_rom_total -1;
	
	function get_next_seed_index (
			index:	in	seed_index_type
		) return seed_index_type;
		
end package seed_table;

package body seed_table is
	
	function get_next_seed_index (
			index:	in	seed_index_type
		) return seed_index_type
	is
	begin
		if index = index'high then
				return 0;
		end if;
		return index + 1;
	end function get_next_seed_index;

end package body seed_table;