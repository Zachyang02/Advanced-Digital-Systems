* run_inverter_nand
.include inverter.cir
.include nand.cir

* subckt for ring_oscillator
.subckt ring_oscillator_2 va in vdd vss

* nand instance
x0 va vb in mid vdd vss nand

* inverter instance
x1 in out vdd vss inverter tplv=65.5n tpwv=216.0n tnln=63.2n tnwm=60.4n tpotv=1.93n tnotv=1.83n
x2 out out2 vdd vss inverter tplv=61.3n tpwv=214.7n tnln=63.4n tnwm=67.8n tpotv=1.92n tnotv=1.83n
x3 out2 out3 vdd vss inverter tplv=58.6n tpwv=212.2n tnln=65.6n tnwm=69.1n tpotv=1.94n tnotv=1.89n
X4 out3 out4 vdd vss inverter tplv=57.2n tpwv=209.6n tnln=62.8n tnwm=67.3n tpotv=1.95n tnotv=1.87n
X5 out4 out5 vdd vss inverter tplv=67.2n tpwv=207.1n tnln=66.8n tnwm=66.6n tpotv=1.94n tnotv=1.86n
X6 out5 out6 vdd vss inverter tplv=66.0n tpwv=212.5n tnln=59.9n tnwm=68.6n tpotv=2.02n tnotv=1.82n
X7 out6 out7 vdd vss inverter tplv=64.5n tpwv=212.2n tnln=59.6n tnwm=66.7n tpotv=1.93n tnotv=1.88n
X8 out7 out8 vdd vss inverter tplv=67.4n tpwv=209.5n tnln=63.9n tnwm=63.9n tpotv=2.0n tnotv=1.86n
X9 out8 out9 vdd vss inverter tplv=61.0n tpwv=219.2n tnln=73.4n tnwm=65.3n tpotv=1.98n tnotv=1.87n
X10 out9 out10 vdd vss inverter tplv=67.3n tpwv=210.0n tnln=59.3n tnwm=63.2n tpotv=2.02n tnotv=1.87n
X11 out10 out11 vdd vss inverter tplv=56.9n tpwv=213.2n tnln=61.1n tnwm=61.8n tpotv=2.0n tnotv=1.86n
X12 out11 vb vdd vss inverter tplv=58.5n tpwv=217.1n tnln=66.4n tnwm=63.3n tpotv=1.96n tnotv=1.83n

.ends ring_oscillator_2