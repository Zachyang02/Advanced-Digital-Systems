library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;





entity top_level is
port();


end entity top_level;



architecture Behavioral of top_level is



begin




end Behavioral;