* run_inverter_nand
.include inverter.cir
.include nand.cir

* subckt for ring_oscillator
.subckt ring_oscillator_7 va in vdd vss

* nand instance
x0 va vb in mid vdd vss nand

* inverter instance
x1 in out vdd vss inverter tplv=68.1n tpwv=213.0n tnln=57.3n tnwm=58.5n tpotv=1.88n tnotv=1.85n
x2 out out2 vdd vss inverter tplv=68.9n tpwv=214.2n tnln=67.8n tnwm=66.2n tpotv=1.91n tnotv=1.82n
x3 out2 out3 vdd vss inverter tplv=64.5n tpwv=221.2n tnln=60.0n tnwm=62.3n tpotv=1.9n tnotv=1.88n
X4 out3 out4 vdd vss inverter tplv=70.5n tpwv=214.4n tnln=59.5n tnwm=64.3n tpotv=1.96n tnotv=1.82n
X5 out4 out5 vdd vss inverter tplv=64.9n tpwv=213.2n tnln=57.9n tnwm=63.0n tpotv=1.95n tnotv=1.83n
X6 out5 out6 vdd vss inverter tplv=63.5n tpwv=210.0n tnln=68.0n tnwm=60.6n tpotv=1.97n tnotv=1.86n
X7 out6 out7 vdd vss inverter tplv=67.3n tpwv=210.2n tnln=69.3n tnwm=69.2n tpotv=1.97n tnotv=1.85n
X8 out7 out8 vdd vss inverter tplv=62.2n tpwv=211.8n tnln=56.6n tnwm=62.5n tpotv=1.94n tnotv=1.8n
X9 out8 out9 vdd vss inverter tplv=61.7n tpwv=217.6n tnln=67.5n tnwm=59.0n tpotv=1.92n tnotv=1.89n
X10 out9 out10 vdd vss inverter tplv=65.4n tpwv=217.2n tnln=64.1n tnwm=67.9n tpotv=1.93n tnotv=1.83n
X11 out10 out11 vdd vss inverter tplv=65.0n tpwv=214.5n tnln=62.8n tnwm=59.7n tpotv=1.97n tnotv=1.84n
X12 out11 vb vdd vss inverter tplv=66.7n tpwv=213.4n tnln=64.9n tnwm=65.5n tpotv=1.95n tnotv=1.84n

.ends ring_oscillator_7