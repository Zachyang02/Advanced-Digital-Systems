* run_inverter_nand
.include inverter.cir
.include nand.cir

* subckt for ring_oscillator
.subckt ring_oscillator_4 va in vdd vss

* nand instance
x0 va vb in mid vdd vss nand

* inverter instance
x1 in out vdd vss inverter tplv=69.0n tpwv=216.7n tnln=58.7n tnwm=60.0n tpotv=1.97n tnotv=1.9n
x2 out out2 vdd vss inverter tplv=69.1n tpwv=218.6n tnln=72.0n tnwm=64.1n tpotv=1.95n tnotv=1.82n
x3 out2 out3 vdd vss inverter tplv=70.9n tpwv=214.4n tnln=59.7n tnwm=65.9n tpotv=1.99n tnotv=1.84n
X4 out3 out4 vdd vss inverter tplv=69.3n tpwv=218.3n tnln=67.9n tnwm=65.0n tpotv=1.95n tnotv=1.85n
X5 out4 out5 vdd vss inverter tplv=63.2n tpwv=214.2n tnln=63.0n tnwm=64.5n tpotv=1.92n tnotv=1.85n
X6 out5 out6 vdd vss inverter tplv=60.4n tpwv=216.5n tnln=72.3n tnwm=69.3n tpotv=1.9n tnotv=1.9n
X7 out6 out7 vdd vss inverter tplv=68.9n tpwv=213.6n tnln=60.1n tnwm=71.0n tpotv=1.92n tnotv=1.84n
X8 out7 out8 vdd vss inverter tplv=64.5n tpwv=216.8n tnln=68.0n tnwm=64.9n tpotv=1.89n tnotv=1.85n
X9 out8 out9 vdd vss inverter tplv=61.7n tpwv=214.1n tnln=66.3n tnwm=64.7n tpotv=1.98n tnotv=1.87n
X10 out9 out10 vdd vss inverter tplv=70.1n tpwv=215.1n tnln=68.0n tnwm=62.6n tpotv=1.95n tnotv=1.85n
X11 out10 out11 vdd vss inverter tplv=71.9n tpwv=208.2n tnln=65.4n tnwm=62.6n tpotv=1.99n tnotv=1.86n
X12 out11 vb vdd vss inverter tplv=66.2n tpwv=215.4n tnln=69.5n tnwm=60.8n tpotv=1.97n tnotv=1.81n

.ends ring_oscillator_4