library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity gen is
    port (

    );
end entity gen;

--In the architecture of the body, you should use a generate statement

architecture mgen of Mandelbrot_gen is
    -- signals
	 
begin

	 
end architecture mgen;