library ads;
use ads.ads_fixed.all;
use ads.ads_complex_pkg.all;

package seed_table is 
	type seed_rom_type is array (natural range<>) of ads_complex;
	constant seed_rom:	seed_rom_type := (
		( re => to_ads_sfixed( 0.00000), im => to_ads_sfixed(-0.00000) ),
			( re => to_ads_sfixed( 0.00748), im => to_ads_sfixed(-0.00748) ),
			( re => to_ads_sfixed( 0.01496), im => to_ads_sfixed(-0.01496) ),
			( re => to_ads_sfixed( 0.02246), im => to_ads_sfixed(-0.02243) ),
			( re => to_ads_sfixed( 0.02996), im => to_ads_sfixed(-0.02990) ),
			( re => to_ads_sfixed( 0.03747), im => to_ads_sfixed(-0.03736) ),
			( re => to_ads_sfixed( 0.04500), im => to_ads_sfixed(-0.04482) ),
			( re => to_ads_sfixed( 0.05255), im => to_ads_sfixed(-0.05226) ),
			( re => to_ads_sfixed( 0.06013), im => to_ads_sfixed(-0.05970) ),
			( re => to_ads_sfixed( 0.06773), im => to_ads_sfixed(-0.06711) ),
			( re => to_ads_sfixed( 0.07536), im => to_ads_sfixed(-0.07452) ),
			( re => to_ads_sfixed( 0.08302), im => to_ads_sfixed(-0.08190) ),
			( re => to_ads_sfixed( 0.09072), im => to_ads_sfixed(-0.08927) ),
			( re => to_ads_sfixed( 0.09847), im => to_ads_sfixed(-0.09661) ),
			( re => to_ads_sfixed( 0.10625), im => to_ads_sfixed(-0.10393) ),
			( re => to_ads_sfixed( 0.11408), im => to_ads_sfixed(-0.11122) ),
			( re => to_ads_sfixed( 0.12197), im => to_ads_sfixed(-0.11849) ),
			( re => to_ads_sfixed( 0.12990), im => to_ads_sfixed(-0.12573) ),
			( re => to_ads_sfixed( 0.13790), im => to_ads_sfixed(-0.13293) ),
			( re => to_ads_sfixed( 0.14595), im => to_ads_sfixed(-0.14010) ),
			( re => to_ads_sfixed( 0.15407), im => to_ads_sfixed(-0.14723) ),
			( re => to_ads_sfixed( 0.16226), im => to_ads_sfixed(-0.15431) ),
			( re => to_ads_sfixed( 0.17051), im => to_ads_sfixed(-0.16136) ),
			( re => to_ads_sfixed( 0.17884), im => to_ads_sfixed(-0.16836) ),
			( re => to_ads_sfixed( 0.18725), im => to_ads_sfixed(-0.17531) ),
			( re => to_ads_sfixed( 0.19573), im => to_ads_sfixed(-0.18220) ),
			( re => to_ads_sfixed( 0.20430), im => to_ads_sfixed(-0.18904) ),
			( re => to_ads_sfixed( 0.21296), im => to_ads_sfixed(-0.19582) ),
			( re => to_ads_sfixed( 0.22171), im => to_ads_sfixed(-0.20254) ),
			( re => to_ads_sfixed( 0.23055), im => to_ads_sfixed(-0.20919) ),
			( re => to_ads_sfixed( 0.23948), im => to_ads_sfixed(-0.21577) ),
			( re => to_ads_sfixed( 0.24852), im => to_ads_sfixed(-0.22227) ),
			( re => to_ads_sfixed( 0.25766), im => to_ads_sfixed(-0.22869) ),
			( re => to_ads_sfixed( 0.26690), im => to_ads_sfixed(-0.23503) ),
			( re => to_ads_sfixed( 0.27625), im => to_ads_sfixed(-0.24128) ),
			( re => to_ads_sfixed( 0.28571), im => to_ads_sfixed(-0.24744) ),
			( re => to_ads_sfixed( 0.29529), im => to_ads_sfixed(-0.25349) ),
			( re => to_ads_sfixed( 0.30498), im => to_ads_sfixed(-0.25944) ),
			( re => to_ads_sfixed( 0.31479), im => to_ads_sfixed(-0.26528) ),
			( re => to_ads_sfixed( 0.32472), im => to_ads_sfixed(-0.27101) ),
			( re => to_ads_sfixed( 0.33478), im => to_ads_sfixed(-0.27661) ),
			( re => to_ads_sfixed( 0.34496), im => to_ads_sfixed(-0.28208) ),
			( re => to_ads_sfixed( 0.35526), im => to_ads_sfixed(-0.28741) ),
			( re => to_ads_sfixed( 0.36570), im => to_ads_sfixed(-0.29261) ),
			( re => to_ads_sfixed( 0.37626), im => to_ads_sfixed(-0.29765) ),
			( re => to_ads_sfixed( 0.38696), im => to_ads_sfixed(-0.30254) ),
			( re => to_ads_sfixed( 0.39779), im => to_ads_sfixed(-0.30726) ),
			( re => to_ads_sfixed( 0.40875), im => to_ads_sfixed(-0.31180) ),
			( re => to_ads_sfixed( 0.41984), im => to_ads_sfixed(-0.31617) ),
			( re => to_ads_sfixed( 0.43107), im => to_ads_sfixed(-0.32035) ),
			( re => to_ads_sfixed( 0.44243), im => to_ads_sfixed(-0.32432) ),
			( re => to_ads_sfixed( 0.45392), im => to_ads_sfixed(-0.32809) ),
			( re => to_ads_sfixed( 0.46554), im => to_ads_sfixed(-0.33164) ),
			( re => to_ads_sfixed( 0.47730), im => to_ads_sfixed(-0.33497) ),
			( re => to_ads_sfixed( 0.48918), im => to_ads_sfixed(-0.33805) ),
			( re => to_ads_sfixed( 0.50119), im => to_ads_sfixed(-0.34089) ),
			( re => to_ads_sfixed( 0.51332), im => to_ads_sfixed(-0.34347) ),
			( re => to_ads_sfixed( 0.52556), im => to_ads_sfixed(-0.34579) ),
			( re => to_ads_sfixed( 0.53793), im => to_ads_sfixed(-0.34782) ),
			( re => to_ads_sfixed( 0.55040), im => to_ads_sfixed(-0.34957) ),
			( re => to_ads_sfixed( 0.56298), im => to_ads_sfixed(-0.35101) ),
			( re => to_ads_sfixed( 0.57566), im => to_ads_sfixed(-0.35214) ),
			( re => to_ads_sfixed( 0.58843), im => to_ads_sfixed(-0.35295) ),
			( re => to_ads_sfixed( 0.60128), im => to_ads_sfixed(-0.35342) ),
			( re => to_ads_sfixed( 0.61421), im => to_ads_sfixed(-0.35355) ),
			( re => to_ads_sfixed( 0.62721), im => to_ads_sfixed(-0.35332) ),
			( re => to_ads_sfixed( 0.64026), im => to_ads_sfixed(-0.35272) ),
			( re => to_ads_sfixed( 0.65336), im => to_ads_sfixed(-0.35174) ),
			( re => to_ads_sfixed( 0.66650), im => to_ads_sfixed(-0.35037) ),
			( re => to_ads_sfixed( 0.67965), im => to_ads_sfixed(-0.34859) ),
			( re => to_ads_sfixed( 0.69282), im => to_ads_sfixed(-0.34641) ),
			( re => to_ads_sfixed( 0.70598), im => to_ads_sfixed(-0.34380) ),
			( re => to_ads_sfixed( 0.71912), im => to_ads_sfixed(-0.34077) ),
			( re => to_ads_sfixed( 0.73222), im => to_ads_sfixed(-0.33729) ),
			( re => to_ads_sfixed( 0.74526), im => to_ads_sfixed(-0.33336) ),
			( re => to_ads_sfixed( 0.75823), im => to_ads_sfixed(-0.32898) ),
			( re => to_ads_sfixed( 0.77110), im => to_ads_sfixed(-0.32414) ),
			( re => to_ads_sfixed( 0.78387), im => to_ads_sfixed(-0.31883) ),
			( re => to_ads_sfixed( 0.79649), im => to_ads_sfixed(-0.31304) ),
			( re => to_ads_sfixed( 0.80897), im => to_ads_sfixed(-0.30678) ),
			( re => to_ads_sfixed( 0.82126), im => to_ads_sfixed(-0.30004) ),
			( re => to_ads_sfixed( 0.83335), im => to_ads_sfixed(-0.29282) ),
			( re => to_ads_sfixed( 0.84521), im => to_ads_sfixed(-0.28511) ),
			( re => to_ads_sfixed( 0.85682), im => to_ads_sfixed(-0.27693) ),
			( re => to_ads_sfixed( 0.86816), im => to_ads_sfixed(-0.26827) ),
			( re => to_ads_sfixed( 0.87919), im => to_ads_sfixed(-0.25915) ),
			( re => to_ads_sfixed( 0.88989), im => to_ads_sfixed(-0.24955) ),
			( re => to_ads_sfixed( 0.90025), im => to_ads_sfixed(-0.23950) ),
			( re => to_ads_sfixed( 0.91022), im => to_ads_sfixed(-0.22900) ),
			( re => to_ads_sfixed( 0.91979), im => to_ads_sfixed(-0.21806) ),
			( re => to_ads_sfixed( 0.92893), im => to_ads_sfixed(-0.20671) ),
			( re => to_ads_sfixed( 0.93762), im => to_ads_sfixed(-0.19494) ),
			( re => to_ads_sfixed( 0.94582), im => to_ads_sfixed(-0.18279) ),
			( re => to_ads_sfixed( 0.95353), im => to_ads_sfixed(-0.17026) ),
			( re => to_ads_sfixed( 0.96071), im => to_ads_sfixed(-0.15738) ),
			( re => to_ads_sfixed( 0.96734), im => to_ads_sfixed(-0.14417) ),
			( re => to_ads_sfixed( 0.97341), im => to_ads_sfixed(-0.13066) ),
			( re => to_ads_sfixed( 0.97889), im => to_ads_sfixed(-0.11687) ),
			( re => to_ads_sfixed( 0.98377), im => to_ads_sfixed(-0.10283) ),
			( re => to_ads_sfixed( 0.98804), im => to_ads_sfixed(-0.08857) ),
			( re => to_ads_sfixed( 0.99167), im => to_ads_sfixed(-0.07411) ),
			( re => to_ads_sfixed( 0.99465), im => to_ads_sfixed(-0.05948) ),
			( re => to_ads_sfixed( 0.99699), im => to_ads_sfixed(-0.04473) ),
			( re => to_ads_sfixed( 0.99866), im => to_ads_sfixed(-0.02988) ),
			( re => to_ads_sfixed( 0.99966), im => to_ads_sfixed(-0.01495) ),
			( re => to_ads_sfixed( 1.00000), im => to_ads_sfixed(-0.00000) ),
			( re => to_ads_sfixed( 0.99966), im => to_ads_sfixed( 0.01495) ),
			( re => to_ads_sfixed( 0.99866), im => to_ads_sfixed( 0.02988) ),
			( re => to_ads_sfixed( 0.99699), im => to_ads_sfixed( 0.04473) ),
			( re => to_ads_sfixed( 0.99465), im => to_ads_sfixed( 0.05948) ),
			( re => to_ads_sfixed( 0.99167), im => to_ads_sfixed( 0.07411) ),
			( re => to_ads_sfixed( 0.98804), im => to_ads_sfixed( 0.08857) ),
			( re => to_ads_sfixed( 0.98377), im => to_ads_sfixed( 0.10283) ),
			( re => to_ads_sfixed( 0.97889), im => to_ads_sfixed( 0.11687) ),
			( re => to_ads_sfixed( 0.97341), im => to_ads_sfixed( 0.13066) ),
			( re => to_ads_sfixed( 0.96734), im => to_ads_sfixed( 0.14417) ),
			( re => to_ads_sfixed( 0.96071), im => to_ads_sfixed( 0.15738) ),
			( re => to_ads_sfixed( 0.95353), im => to_ads_sfixed( 0.17026) ),
			( re => to_ads_sfixed( 0.94582), im => to_ads_sfixed( 0.18279) ),
			( re => to_ads_sfixed( 0.93762), im => to_ads_sfixed( 0.19494) ),
			( re => to_ads_sfixed( 0.92893), im => to_ads_sfixed( 0.20671) ),
			( re => to_ads_sfixed( 0.91979), im => to_ads_sfixed( 0.21806) ),
			( re => to_ads_sfixed( 0.91022), im => to_ads_sfixed( 0.22900) ),
			( re => to_ads_sfixed( 0.90025), im => to_ads_sfixed( 0.23950) ),
			( re => to_ads_sfixed( 0.88989), im => to_ads_sfixed( 0.24955) ),
			( re => to_ads_sfixed( 0.87919), im => to_ads_sfixed( 0.25915) ),
			( re => to_ads_sfixed( 0.86816), im => to_ads_sfixed( 0.26827) ),
			( re => to_ads_sfixed( 0.85682), im => to_ads_sfixed( 0.27693) ),
			( re => to_ads_sfixed( 0.84521), im => to_ads_sfixed( 0.28511) ),
			( re => to_ads_sfixed( 0.83335), im => to_ads_sfixed( 0.29282) ),
			( re => to_ads_sfixed( 0.82126), im => to_ads_sfixed( 0.30004) ),
			( re => to_ads_sfixed( 0.80897), im => to_ads_sfixed( 0.30678) ),
			( re => to_ads_sfixed( 0.79649), im => to_ads_sfixed( 0.31304) ),
			( re => to_ads_sfixed( 0.78387), im => to_ads_sfixed( 0.31883) ),
			( re => to_ads_sfixed( 0.77110), im => to_ads_sfixed( 0.32414) ),
			( re => to_ads_sfixed( 0.75823), im => to_ads_sfixed( 0.32898) ),
			( re => to_ads_sfixed( 0.74526), im => to_ads_sfixed( 0.33336) ),
			( re => to_ads_sfixed( 0.73222), im => to_ads_sfixed( 0.33729) ),
			( re => to_ads_sfixed( 0.71912), im => to_ads_sfixed( 0.34077) ),
			( re => to_ads_sfixed( 0.70598), im => to_ads_sfixed( 0.34380) ),
			( re => to_ads_sfixed( 0.69282), im => to_ads_sfixed( 0.34641) ),
			( re => to_ads_sfixed( 0.67965), im => to_ads_sfixed( 0.34859) ),
			( re => to_ads_sfixed( 0.66650), im => to_ads_sfixed( 0.35037) ),
			( re => to_ads_sfixed( 0.65336), im => to_ads_sfixed( 0.35174) ),
			( re => to_ads_sfixed( 0.64026), im => to_ads_sfixed( 0.35272) ),
			( re => to_ads_sfixed( 0.62721), im => to_ads_sfixed( 0.35332) ),
			( re => to_ads_sfixed( 0.61421), im => to_ads_sfixed( 0.35355) ),
			( re => to_ads_sfixed( 0.60128), im => to_ads_sfixed( 0.35342) ),
			( re => to_ads_sfixed( 0.58843), im => to_ads_sfixed( 0.35295) ),
			( re => to_ads_sfixed( 0.57566), im => to_ads_sfixed( 0.35214) ),
			( re => to_ads_sfixed( 0.56298), im => to_ads_sfixed( 0.35101) ),
			( re => to_ads_sfixed( 0.55040), im => to_ads_sfixed( 0.34957) ),
			( re => to_ads_sfixed( 0.53793), im => to_ads_sfixed( 0.34782) ),
			( re => to_ads_sfixed( 0.52556), im => to_ads_sfixed( 0.34579) ),
			( re => to_ads_sfixed( 0.51332), im => to_ads_sfixed( 0.34347) ),
			( re => to_ads_sfixed( 0.50119), im => to_ads_sfixed( 0.34089) ),
			( re => to_ads_sfixed( 0.48918), im => to_ads_sfixed( 0.33805) ),
			( re => to_ads_sfixed( 0.47730), im => to_ads_sfixed( 0.33497) ),
			( re => to_ads_sfixed( 0.46554), im => to_ads_sfixed( 0.33164) ),
			( re => to_ads_sfixed( 0.45392), im => to_ads_sfixed( 0.32809) ),
			( re => to_ads_sfixed( 0.44243), im => to_ads_sfixed( 0.32432) ),
			( re => to_ads_sfixed( 0.43107), im => to_ads_sfixed( 0.32035) ),
			( re => to_ads_sfixed( 0.41984), im => to_ads_sfixed( 0.31617) ),
			( re => to_ads_sfixed( 0.40875), im => to_ads_sfixed( 0.31180) ),
			( re => to_ads_sfixed( 0.39779), im => to_ads_sfixed( 0.30726) ),
			( re => to_ads_sfixed( 0.38696), im => to_ads_sfixed( 0.30254) ),
			( re => to_ads_sfixed( 0.37626), im => to_ads_sfixed( 0.29765) ),
			( re => to_ads_sfixed( 0.36570), im => to_ads_sfixed( 0.29261) ),
			( re => to_ads_sfixed( 0.35526), im => to_ads_sfixed( 0.28741) ),
			( re => to_ads_sfixed( 0.34496), im => to_ads_sfixed( 0.28208) ),
			( re => to_ads_sfixed( 0.33478), im => to_ads_sfixed( 0.27661) ),
			( re => to_ads_sfixed( 0.32472), im => to_ads_sfixed( 0.27101) ),
			( re => to_ads_sfixed( 0.31479), im => to_ads_sfixed( 0.26528) ),
			( re => to_ads_sfixed( 0.30498), im => to_ads_sfixed( 0.25944) ),
			( re => to_ads_sfixed( 0.29529), im => to_ads_sfixed( 0.25349) ),
			( re => to_ads_sfixed( 0.28571), im => to_ads_sfixed( 0.24744) ),
			( re => to_ads_sfixed( 0.27625), im => to_ads_sfixed( 0.24128) ),
			( re => to_ads_sfixed( 0.26690), im => to_ads_sfixed( 0.23503) ),
			( re => to_ads_sfixed( 0.25766), im => to_ads_sfixed( 0.22869) ),
			( re => to_ads_sfixed( 0.24852), im => to_ads_sfixed( 0.22227) ),
			( re => to_ads_sfixed( 0.23948), im => to_ads_sfixed( 0.21577) ),
			( re => to_ads_sfixed( 0.23055), im => to_ads_sfixed( 0.20919) ),
			( re => to_ads_sfixed( 0.22171), im => to_ads_sfixed( 0.20254) ),
			( re => to_ads_sfixed( 0.21296), im => to_ads_sfixed( 0.19582) ),
			( re => to_ads_sfixed( 0.20430), im => to_ads_sfixed( 0.18904) ),
			( re => to_ads_sfixed( 0.19573), im => to_ads_sfixed( 0.18220) ),
			( re => to_ads_sfixed( 0.18725), im => to_ads_sfixed( 0.17531) ),
			( re => to_ads_sfixed( 0.17884), im => to_ads_sfixed( 0.16836) ),
			( re => to_ads_sfixed( 0.17051), im => to_ads_sfixed( 0.16136) ),
			( re => to_ads_sfixed( 0.16226), im => to_ads_sfixed( 0.15431) ),
			( re => to_ads_sfixed( 0.15407), im => to_ads_sfixed( 0.14723) ),
			( re => to_ads_sfixed( 0.14595), im => to_ads_sfixed( 0.14010) ),
			( re => to_ads_sfixed( 0.13790), im => to_ads_sfixed( 0.13293) ),
			( re => to_ads_sfixed( 0.12990), im => to_ads_sfixed( 0.12573) ),
			( re => to_ads_sfixed( 0.12197), im => to_ads_sfixed( 0.11849) ),
			( re => to_ads_sfixed( 0.11408), im => to_ads_sfixed( 0.11122) ),
			( re => to_ads_sfixed( 0.10625), im => to_ads_sfixed( 0.10393) ),
			( re => to_ads_sfixed( 0.09847), im => to_ads_sfixed( 0.09661) ),
			( re => to_ads_sfixed( 0.09072), im => to_ads_sfixed( 0.08927) ),
			( re => to_ads_sfixed( 0.08302), im => to_ads_sfixed( 0.08190) ),
			( re => to_ads_sfixed( 0.07536), im => to_ads_sfixed( 0.07452) ),
			( re => to_ads_sfixed( 0.06773), im => to_ads_sfixed( 0.06711) ),
			( re => to_ads_sfixed( 0.06013), im => to_ads_sfixed( 0.05970) ),
			( re => to_ads_sfixed( 0.05255), im => to_ads_sfixed( 0.05226) ),
			( re => to_ads_sfixed( 0.04500), im => to_ads_sfixed( 0.04482) ),
			( re => to_ads_sfixed( 0.03747), im => to_ads_sfixed( 0.03736) ),
			( re => to_ads_sfixed( 0.02996), im => to_ads_sfixed( 0.02990) ),
			( re => to_ads_sfixed( 0.02246), im => to_ads_sfixed( 0.02243) ),
			( re => to_ads_sfixed( 0.01496), im => to_ads_sfixed( 0.01496) ),
			( re => to_ads_sfixed( 0.00748), im => to_ads_sfixed( 0.00748) ),
			( re => to_ads_sfixed( 0.00000), im => to_ads_sfixed( 0.00000) ),
			( re => to_ads_sfixed(-0.00748), im => to_ads_sfixed(-0.00748) ),
			( re => to_ads_sfixed(-0.01496), im => to_ads_sfixed(-0.01496) ),
			( re => to_ads_sfixed(-0.02246), im => to_ads_sfixed(-0.02243) ),
			( re => to_ads_sfixed(-0.02996), im => to_ads_sfixed(-0.02990) ),
			( re => to_ads_sfixed(-0.03747), im => to_ads_sfixed(-0.03736) ),
			( re => to_ads_sfixed(-0.04500), im => to_ads_sfixed(-0.04482) ),
			( re => to_ads_sfixed(-0.05255), im => to_ads_sfixed(-0.05226) ),
			( re => to_ads_sfixed(-0.06013), im => to_ads_sfixed(-0.05970) ),
			( re => to_ads_sfixed(-0.06773), im => to_ads_sfixed(-0.06711) ),
			( re => to_ads_sfixed(-0.07536), im => to_ads_sfixed(-0.07452) ),
			( re => to_ads_sfixed(-0.08302), im => to_ads_sfixed(-0.08190) ),
			( re => to_ads_sfixed(-0.09072), im => to_ads_sfixed(-0.08927) ),
			( re => to_ads_sfixed(-0.09847), im => to_ads_sfixed(-0.09661) ),
			( re => to_ads_sfixed(-0.10625), im => to_ads_sfixed(-0.10393) ),
			( re => to_ads_sfixed(-0.11408), im => to_ads_sfixed(-0.11122) ),
			( re => to_ads_sfixed(-0.12197), im => to_ads_sfixed(-0.11849) ),
			( re => to_ads_sfixed(-0.12990), im => to_ads_sfixed(-0.12573) ),
			( re => to_ads_sfixed(-0.13790), im => to_ads_sfixed(-0.13293) ),
			( re => to_ads_sfixed(-0.14595), im => to_ads_sfixed(-0.14010) ),
			( re => to_ads_sfixed(-0.15407), im => to_ads_sfixed(-0.14723) ),
			( re => to_ads_sfixed(-0.16226), im => to_ads_sfixed(-0.15431) ),
			( re => to_ads_sfixed(-0.17051), im => to_ads_sfixed(-0.16136) ),
			( re => to_ads_sfixed(-0.17884), im => to_ads_sfixed(-0.16836) ),
			( re => to_ads_sfixed(-0.18725), im => to_ads_sfixed(-0.17531) ),
			( re => to_ads_sfixed(-0.19573), im => to_ads_sfixed(-0.18220) ),
			( re => to_ads_sfixed(-0.20430), im => to_ads_sfixed(-0.18904) ),
			( re => to_ads_sfixed(-0.21296), im => to_ads_sfixed(-0.19582) ),
			( re => to_ads_sfixed(-0.22171), im => to_ads_sfixed(-0.20254) ),
			( re => to_ads_sfixed(-0.23055), im => to_ads_sfixed(-0.20919) ),
			( re => to_ads_sfixed(-0.23948), im => to_ads_sfixed(-0.21577) ),
			( re => to_ads_sfixed(-0.24852), im => to_ads_sfixed(-0.22227) ),
			( re => to_ads_sfixed(-0.25766), im => to_ads_sfixed(-0.22869) ),
			( re => to_ads_sfixed(-0.26690), im => to_ads_sfixed(-0.23503) ),
			( re => to_ads_sfixed(-0.27625), im => to_ads_sfixed(-0.24128) ),
			( re => to_ads_sfixed(-0.28571), im => to_ads_sfixed(-0.24744) ),
			( re => to_ads_sfixed(-0.29529), im => to_ads_sfixed(-0.25349) ),
			( re => to_ads_sfixed(-0.30498), im => to_ads_sfixed(-0.25944) ),
			( re => to_ads_sfixed(-0.31479), im => to_ads_sfixed(-0.26528) ),
			( re => to_ads_sfixed(-0.32472), im => to_ads_sfixed(-0.27101) ),
			( re => to_ads_sfixed(-0.33478), im => to_ads_sfixed(-0.27661) ),
			( re => to_ads_sfixed(-0.34496), im => to_ads_sfixed(-0.28208) ),
			( re => to_ads_sfixed(-0.35526), im => to_ads_sfixed(-0.28741) ),
			( re => to_ads_sfixed(-0.36570), im => to_ads_sfixed(-0.29261) ),
			( re => to_ads_sfixed(-0.37626), im => to_ads_sfixed(-0.29765) ),
			( re => to_ads_sfixed(-0.38696), im => to_ads_sfixed(-0.30254) ),
			( re => to_ads_sfixed(-0.39779), im => to_ads_sfixed(-0.30726) ),
			( re => to_ads_sfixed(-0.40875), im => to_ads_sfixed(-0.31180) ),
			( re => to_ads_sfixed(-0.41984), im => to_ads_sfixed(-0.31617) ),
			( re => to_ads_sfixed(-0.43107), im => to_ads_sfixed(-0.32035) ),
			( re => to_ads_sfixed(-0.44243), im => to_ads_sfixed(-0.32432) ),
			( re => to_ads_sfixed(-0.45392), im => to_ads_sfixed(-0.32809) ),
			( re => to_ads_sfixed(-0.46554), im => to_ads_sfixed(-0.33164) ),
			( re => to_ads_sfixed(-0.47730), im => to_ads_sfixed(-0.33497) ),
			( re => to_ads_sfixed(-0.48918), im => to_ads_sfixed(-0.33805) ),
			( re => to_ads_sfixed(-0.50119), im => to_ads_sfixed(-0.34089) ),
			( re => to_ads_sfixed(-0.51332), im => to_ads_sfixed(-0.34347) ),
			( re => to_ads_sfixed(-0.52556), im => to_ads_sfixed(-0.34579) ),
			( re => to_ads_sfixed(-0.53793), im => to_ads_sfixed(-0.34782) ),
			( re => to_ads_sfixed(-0.55040), im => to_ads_sfixed(-0.34957) ),
			( re => to_ads_sfixed(-0.56298), im => to_ads_sfixed(-0.35101) ),
			( re => to_ads_sfixed(-0.57566), im => to_ads_sfixed(-0.35214) ),
			( re => to_ads_sfixed(-0.58843), im => to_ads_sfixed(-0.35295) ),
			( re => to_ads_sfixed(-0.60128), im => to_ads_sfixed(-0.35342) ),
			( re => to_ads_sfixed(-0.61421), im => to_ads_sfixed(-0.35355) ),
			( re => to_ads_sfixed(-0.62721), im => to_ads_sfixed(-0.35332) ),
			( re => to_ads_sfixed(-0.64026), im => to_ads_sfixed(-0.35272) ),
			( re => to_ads_sfixed(-0.65336), im => to_ads_sfixed(-0.35174) ),
			( re => to_ads_sfixed(-0.66650), im => to_ads_sfixed(-0.35037) ),
			( re => to_ads_sfixed(-0.67965), im => to_ads_sfixed(-0.34859) ),
			( re => to_ads_sfixed(-0.69282), im => to_ads_sfixed(-0.34641) ),
			( re => to_ads_sfixed(-0.70598), im => to_ads_sfixed(-0.34380) ),
			( re => to_ads_sfixed(-0.71912), im => to_ads_sfixed(-0.34077) ),
			( re => to_ads_sfixed(-0.73222), im => to_ads_sfixed(-0.33729) ),
			( re => to_ads_sfixed(-0.74526), im => to_ads_sfixed(-0.33336) ),
			( re => to_ads_sfixed(-0.75823), im => to_ads_sfixed(-0.32898) ),
			( re => to_ads_sfixed(-0.77110), im => to_ads_sfixed(-0.32414) ),
			( re => to_ads_sfixed(-0.78387), im => to_ads_sfixed(-0.31883) ),
			( re => to_ads_sfixed(-0.79649), im => to_ads_sfixed(-0.31304) ),
			( re => to_ads_sfixed(-0.80897), im => to_ads_sfixed(-0.30678) ),
			( re => to_ads_sfixed(-0.82126), im => to_ads_sfixed(-0.30004) ),
			( re => to_ads_sfixed(-0.83335), im => to_ads_sfixed(-0.29282) ),
			( re => to_ads_sfixed(-0.84521), im => to_ads_sfixed(-0.28511) ),
			( re => to_ads_sfixed(-0.85682), im => to_ads_sfixed(-0.27693) ),
			( re => to_ads_sfixed(-0.86816), im => to_ads_sfixed(-0.26827) ),
			( re => to_ads_sfixed(-0.87919), im => to_ads_sfixed(-0.25915) ),
			( re => to_ads_sfixed(-0.88989), im => to_ads_sfixed(-0.24955) ),
			( re => to_ads_sfixed(-0.90025), im => to_ads_sfixed(-0.23950) ),
			( re => to_ads_sfixed(-0.91022), im => to_ads_sfixed(-0.22900) ),
			( re => to_ads_sfixed(-0.91979), im => to_ads_sfixed(-0.21806) ),
			( re => to_ads_sfixed(-0.92893), im => to_ads_sfixed(-0.20671) ),
			( re => to_ads_sfixed(-0.93762), im => to_ads_sfixed(-0.19494) ),
			( re => to_ads_sfixed(-0.94582), im => to_ads_sfixed(-0.18279) ),
			( re => to_ads_sfixed(-0.95353), im => to_ads_sfixed(-0.17026) ),
			( re => to_ads_sfixed(-0.96071), im => to_ads_sfixed(-0.15738) ),
			( re => to_ads_sfixed(-0.96734), im => to_ads_sfixed(-0.14417) ),
			( re => to_ads_sfixed(-0.97341), im => to_ads_sfixed(-0.13066) ),
			( re => to_ads_sfixed(-0.97889), im => to_ads_sfixed(-0.11687) ),
			( re => to_ads_sfixed(-0.98377), im => to_ads_sfixed(-0.10283) ),
			( re => to_ads_sfixed(-0.98804), im => to_ads_sfixed(-0.08857) ),
			( re => to_ads_sfixed(-0.99167), im => to_ads_sfixed(-0.07411) ),
			( re => to_ads_sfixed(-0.99465), im => to_ads_sfixed(-0.05948) ),
			( re => to_ads_sfixed(-0.99699), im => to_ads_sfixed(-0.04473) ),
			( re => to_ads_sfixed(-0.99866), im => to_ads_sfixed(-0.02988) ),
			( re => to_ads_sfixed(-0.99966), im => to_ads_sfixed(-0.01495) ),
			( re => to_ads_sfixed(-1.00000), im => to_ads_sfixed( 0.00000) ),
			( re => to_ads_sfixed(-0.99966), im => to_ads_sfixed( 0.01495) ),
			( re => to_ads_sfixed(-0.99866), im => to_ads_sfixed( 0.02988) ),
			( re => to_ads_sfixed(-0.99699), im => to_ads_sfixed( 0.04473) ),
			( re => to_ads_sfixed(-0.99465), im => to_ads_sfixed( 0.05948) ),
			( re => to_ads_sfixed(-0.99167), im => to_ads_sfixed( 0.07411) ),
			( re => to_ads_sfixed(-0.98804), im => to_ads_sfixed( 0.08857) ),
			( re => to_ads_sfixed(-0.98377), im => to_ads_sfixed( 0.10283) ),
			( re => to_ads_sfixed(-0.97889), im => to_ads_sfixed( 0.11687) ),
			( re => to_ads_sfixed(-0.97341), im => to_ads_sfixed( 0.13066) ),
			( re => to_ads_sfixed(-0.96734), im => to_ads_sfixed( 0.14417) ),
			( re => to_ads_sfixed(-0.96071), im => to_ads_sfixed( 0.15738) ),
			( re => to_ads_sfixed(-0.95353), im => to_ads_sfixed( 0.17026) ),
			( re => to_ads_sfixed(-0.94582), im => to_ads_sfixed( 0.18279) ),
			( re => to_ads_sfixed(-0.93762), im => to_ads_sfixed( 0.19494) ),
			( re => to_ads_sfixed(-0.92893), im => to_ads_sfixed( 0.20671) ),
			( re => to_ads_sfixed(-0.91979), im => to_ads_sfixed( 0.21806) ),
			( re => to_ads_sfixed(-0.91022), im => to_ads_sfixed( 0.22900) ),
			( re => to_ads_sfixed(-0.90025), im => to_ads_sfixed( 0.23950) ),
			( re => to_ads_sfixed(-0.88989), im => to_ads_sfixed( 0.24955) ),
			( re => to_ads_sfixed(-0.87919), im => to_ads_sfixed( 0.25915) ),
			( re => to_ads_sfixed(-0.86816), im => to_ads_sfixed( 0.26827) ),
			( re => to_ads_sfixed(-0.85682), im => to_ads_sfixed( 0.27693) ),
			( re => to_ads_sfixed(-0.84521), im => to_ads_sfixed( 0.28511) ),
			( re => to_ads_sfixed(-0.83335), im => to_ads_sfixed( 0.29282) ),
			( re => to_ads_sfixed(-0.82126), im => to_ads_sfixed( 0.30004) ),
			( re => to_ads_sfixed(-0.80897), im => to_ads_sfixed( 0.30678) ),
			( re => to_ads_sfixed(-0.79649), im => to_ads_sfixed( 0.31304) ),
			( re => to_ads_sfixed(-0.78387), im => to_ads_sfixed( 0.31883) ),
			( re => to_ads_sfixed(-0.77110), im => to_ads_sfixed( 0.32414) ),
			( re => to_ads_sfixed(-0.75823), im => to_ads_sfixed( 0.32898) ),
			( re => to_ads_sfixed(-0.74526), im => to_ads_sfixed( 0.33336) ),
			( re => to_ads_sfixed(-0.73222), im => to_ads_sfixed( 0.33729) ),
			( re => to_ads_sfixed(-0.71912), im => to_ads_sfixed( 0.34077) ),
			( re => to_ads_sfixed(-0.70598), im => to_ads_sfixed( 0.34380) ),
			( re => to_ads_sfixed(-0.69282), im => to_ads_sfixed( 0.34641) ),
			( re => to_ads_sfixed(-0.67965), im => to_ads_sfixed( 0.34859) ),
			( re => to_ads_sfixed(-0.66650), im => to_ads_sfixed( 0.35037) ),
			( re => to_ads_sfixed(-0.65336), im => to_ads_sfixed( 0.35174) ),
			( re => to_ads_sfixed(-0.64026), im => to_ads_sfixed( 0.35272) ),
			( re => to_ads_sfixed(-0.62721), im => to_ads_sfixed( 0.35332) ),
			( re => to_ads_sfixed(-0.61421), im => to_ads_sfixed( 0.35355) ),
			( re => to_ads_sfixed(-0.60128), im => to_ads_sfixed( 0.35342) ),
			( re => to_ads_sfixed(-0.58843), im => to_ads_sfixed( 0.35295) ),
			( re => to_ads_sfixed(-0.57566), im => to_ads_sfixed( 0.35214) ),
			( re => to_ads_sfixed(-0.56298), im => to_ads_sfixed( 0.35101) ),
			( re => to_ads_sfixed(-0.55040), im => to_ads_sfixed( 0.34957) ),
			( re => to_ads_sfixed(-0.53793), im => to_ads_sfixed( 0.34782) ),
			( re => to_ads_sfixed(-0.52556), im => to_ads_sfixed( 0.34579) ),
			( re => to_ads_sfixed(-0.51332), im => to_ads_sfixed( 0.34347) ),
			( re => to_ads_sfixed(-0.50119), im => to_ads_sfixed( 0.34089) ),
			( re => to_ads_sfixed(-0.48918), im => to_ads_sfixed( 0.33805) ),
			( re => to_ads_sfixed(-0.47730), im => to_ads_sfixed( 0.33497) ),
			( re => to_ads_sfixed(-0.46554), im => to_ads_sfixed( 0.33164) ),
			( re => to_ads_sfixed(-0.45392), im => to_ads_sfixed( 0.32809) ),
			( re => to_ads_sfixed(-0.44243), im => to_ads_sfixed( 0.32432) ),
			( re => to_ads_sfixed(-0.43107), im => to_ads_sfixed( 0.32035) ),
			( re => to_ads_sfixed(-0.41984), im => to_ads_sfixed( 0.31617) ),
			( re => to_ads_sfixed(-0.40875), im => to_ads_sfixed( 0.31180) ),
			( re => to_ads_sfixed(-0.39779), im => to_ads_sfixed( 0.30726) ),
			( re => to_ads_sfixed(-0.38696), im => to_ads_sfixed( 0.30254) ),
			( re => to_ads_sfixed(-0.37626), im => to_ads_sfixed( 0.29765) ),
			( re => to_ads_sfixed(-0.36570), im => to_ads_sfixed( 0.29261) ),
			( re => to_ads_sfixed(-0.35526), im => to_ads_sfixed( 0.28741) ),
			( re => to_ads_sfixed(-0.34496), im => to_ads_sfixed( 0.28208) ),
			( re => to_ads_sfixed(-0.33478), im => to_ads_sfixed( 0.27661) ),
			( re => to_ads_sfixed(-0.32472), im => to_ads_sfixed( 0.27101) ),
			( re => to_ads_sfixed(-0.31479), im => to_ads_sfixed( 0.26528) ),
			( re => to_ads_sfixed(-0.30498), im => to_ads_sfixed( 0.25944) ),
			( re => to_ads_sfixed(-0.29529), im => to_ads_sfixed( 0.25349) ),
			( re => to_ads_sfixed(-0.28571), im => to_ads_sfixed( 0.24744) ),
			( re => to_ads_sfixed(-0.27625), im => to_ads_sfixed( 0.24128) ),
			( re => to_ads_sfixed(-0.26690), im => to_ads_sfixed( 0.23503) ),
			( re => to_ads_sfixed(-0.25766), im => to_ads_sfixed( 0.22869) ),
			( re => to_ads_sfixed(-0.24852), im => to_ads_sfixed( 0.22227) ),
			( re => to_ads_sfixed(-0.23948), im => to_ads_sfixed( 0.21577) ),
			( re => to_ads_sfixed(-0.23055), im => to_ads_sfixed( 0.20919) ),
			( re => to_ads_sfixed(-0.22171), im => to_ads_sfixed( 0.20254) ),
			( re => to_ads_sfixed(-0.21296), im => to_ads_sfixed( 0.19582) ),
			( re => to_ads_sfixed(-0.20430), im => to_ads_sfixed( 0.18904) ),
			( re => to_ads_sfixed(-0.19573), im => to_ads_sfixed( 0.18220) ),
			( re => to_ads_sfixed(-0.18725), im => to_ads_sfixed( 0.17531) ),
			( re => to_ads_sfixed(-0.17884), im => to_ads_sfixed( 0.16836) ),
			( re => to_ads_sfixed(-0.17051), im => to_ads_sfixed( 0.16136) ),
			( re => to_ads_sfixed(-0.16226), im => to_ads_sfixed( 0.15431) ),
			( re => to_ads_sfixed(-0.15407), im => to_ads_sfixed( 0.14723) ),
			( re => to_ads_sfixed(-0.14595), im => to_ads_sfixed( 0.14010) ),
			( re => to_ads_sfixed(-0.13790), im => to_ads_sfixed( 0.13293) ),
			( re => to_ads_sfixed(-0.12990), im => to_ads_sfixed( 0.12573) ),
			( re => to_ads_sfixed(-0.12197), im => to_ads_sfixed( 0.11849) ),
			( re => to_ads_sfixed(-0.11408), im => to_ads_sfixed( 0.11122) ),
			( re => to_ads_sfixed(-0.10625), im => to_ads_sfixed( 0.10393) ),
			( re => to_ads_sfixed(-0.09847), im => to_ads_sfixed( 0.09661) ),
			( re => to_ads_sfixed(-0.09072), im => to_ads_sfixed( 0.08927) ),
			( re => to_ads_sfixed(-0.08302), im => to_ads_sfixed( 0.08190) ),
			( re => to_ads_sfixed(-0.07536), im => to_ads_sfixed( 0.07452) ),
			( re => to_ads_sfixed(-0.06773), im => to_ads_sfixed( 0.06711) ),
			( re => to_ads_sfixed(-0.06013), im => to_ads_sfixed( 0.05970) ),
			( re => to_ads_sfixed(-0.05255), im => to_ads_sfixed( 0.05226) ),
			( re => to_ads_sfixed(-0.04500), im => to_ads_sfixed( 0.04482) ),
			( re => to_ads_sfixed(-0.03747), im => to_ads_sfixed( 0.03736) ),
			( re => to_ads_sfixed(-0.02996), im => to_ads_sfixed( 0.02990) ),
			( re => to_ads_sfixed(-0.02246), im => to_ads_sfixed( 0.02243) ),
			( re => to_ads_sfixed(-0.01496), im => to_ads_sfixed( 0.01496) ),
			( re => to_ads_sfixed(-0.00748), im => to_ads_sfixed( 0.00748) )
	);
	
	
	constant seed_rom_total: natural := seed_rom'length;
	
	
	subtype seed_index_type is natural range 0 to seed_rom_total -1;
	
	function get_next_seed_index (
			index:	in	seed_index_type
		) return seed_index_type;
		
end package seed_table;

package body seed_table is
	
	function get_next_seed_index (
			index:	in	seed_index_type
		) return seed_index_type
	is
	begin
		if index = index'high then
				return 0;
		end if;
		return index + 1;
	end function get_next_seed_index;

end package body seed_table;